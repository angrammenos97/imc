`define SOC_MEM_MAP_PEC_START_ADDR  32'h1A40_0000
`define SOC_MEM_MAP_PEC_END_ADDR    32'h1A40_1000
