`include "register_interface/typedef.svh"
`include "register_interface/assign.svh"

module pec_axi_to_ip
    import pec_reg_pkg::pec_reg2hw_t;
    import pec_reg_pkg::pec_hw2reg_t;
#(
    parameter int unsigned AXI_ADDR_WIDTH   = 32,
    parameter int unsigned AXI_DATA_WIDTH   = 32,
    parameter int unsigned AXI_ID_WIDTH     = -1,
    parameter int unsigned AXI_USER_WIDTH   = -1
) (
    input logic         clk_i,
    input logic         rst_ni,
    input logic         test_mode_i,
    input pec_hw2reg_t  ip_to_reg_file_i,
    AXI_BUS.Slave       slv,
    output pec_reg2hw_t reg_file_to_ip_o
);

    REG_BUS #(
        .ADDR_WIDTH(AXI_ADDR_WIDTH), 
        .DATA_WIDTH(AXI_DATA_WIDTH)
    ) axi_to_reg_file (
        .clk_i(clk_i)
    );

    //Convert the REG_BUS interface to the struct signals used by the autogenerated interface
    typedef logic [AXI_DATA_WIDTH-1:0] data_t;
    typedef logic [AXI_ADDR_WIDTH-1:0] addr_t;
    typedef logic [AXI_DATA_WIDTH/8-1:0] strb_t;
    `REG_BUS_TYPEDEF_REQ(reg_req_t, addr_t, data_t, strb_t)
    `REG_BUS_TYPEDEF_RSP(reg_rsp_t, data_t)
    reg_req_t to_reg_file_req;
    reg_rsp_t from_reg_file_rsp;
    `REG_BUS_ASSIGN_TO_REQ(to_reg_file_req, axi_to_reg_file)
    `REG_BUS_ASSIGN_FROM_RSP(axi_to_reg_file, from_reg_file_rsp)

    axi_to_reg_intf #(
        .ADDR_WIDTH (AXI_ADDR_WIDTH),
        .DATA_WIDTH (AXI_DATA_WIDTH),
        .ID_WIDTH   (AXI_ID_WIDTH),
        .USER_WIDTH (AXI_USER_WIDTH),
        .DECOUPLE_W (0)
    ) axi_to_reg_intf_i (
        .clk_i      (clk_i),
        .rst_ni     (rst_ni),
        .testmode_i (test_mode_i),
        .in         (slv),
        .reg_o      (axi_to_reg_file)
    );

    pec_reg_top #(
        .reg_req_t(reg_req_t),
        .reg_rsp_t(reg_rsp_t)
    ) pec_reg_top_i (
        .clk_i      (clk_i),
        .rst_ni     (rst_ni),
        .reg_req_i  (to_reg_file_req),
        .reg_rsp_o  (from_reg_file_rsp),
        .reg2hw     (reg_file_to_ip_o),
        .hw2reg     (ip_to_reg_file_i),
        .devmode_i  (1'b1)
    );

endmodule